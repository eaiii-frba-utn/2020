* C:\Audio\TubeShar\Pent_P.sch

* Schematics Version 6.3 - April 1996
* Sun Sep 02 12:29:32 2001


** Analysis setup **
.DC LIN V_VP 0 600 5 
.STEP LIN V_VG1 0 -50 -10 


* From [SCHEMATICS NETLIST] section of msim.ini:
.lib C:\AUDIO\TubeShar\TUBE.LIB
.lib nom.lib

.INC "Pent_P.net"
.INC "Pent_P.als"


.probe


.END
